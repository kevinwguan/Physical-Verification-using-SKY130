** sch_path: /home/kevin/Documents/Day1/inverter/xschem/inverter_tb.sch
**.subckt inverter_tb in out
*.opin in
*.opin out
x1 net1 in out GND inverter
V1 in GND PWL(0 0 500n 0 1000n 1.8 1500n 1.8)
.save i(v1)
V2 net1 GND 1.8
.save i(v2)
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 1n 2u
plot v(in) v(out)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/kevin/Documents/Day1/inverter/xschem/inverter.sym
** sch_path: /home/kevin/Documents/Day1/inverter/xschem/inverter.sch
.subckt inverter vdd in out vss
*.ipin in
*.iopin vdd
*.iopin vss
*.opin out
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=13.5 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd VDD sky130_fd_pr__pfet_01v8 L=0.18 W=9 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.save all
.GLOBAL GND
.end
